// The environment is a container object simply to hold all verification 
// components together. This environment can then be reused later and all
// components in it would be automatically connected and available for use
// This is an environment without a generator.
class env;
    driver 			d0; 		// Driver to design
    monitor 			m0; 		// Monitor from design
    scoreboard 		s0; 		// Scoreboard connected to monitor
    mailbox 			scb_mbx; 	// Top level mailbox for SCB <-> MON 
    virtual reg_if 	vif; 		// Virtual interface handle

    // Instantiate all testbench components
    function new();
        d0 = new;
        m0 = new;
        s0 = new;
        scb_mbx = new();
    endfunction

    // Assign handles and start all components so that 
    // they all become active and wait for transactions to be
    // available
    virtual task run();
        d0.vif = vif;
        m0.vif = vif;
        m0.scb_mbx = scb_mbx;
        s0.scb_mbx = scb_mbx;
        
        fork
            s0.run();
            d0.run();
            m0.run();
        join_any
    endtask
    endclass

    // Sometimes we simply need to generate N random transactions to random
    // locations so a generator would be useful to do just that. In this case
    // loop determines how many transactions need to be sent
    class generator;
    int 	loop = 10;
    event drv_done;
    mailbox drv_mbx;

    task run();
        for (int i = 0; i < loop; i++) begin
        reg_item item = new;
        item.randomize();
        $display ("T=%0t [Generator] Loop:%0d/%0d create next item", $time, i+1, loop);
        drv_mbx.put(item);
        $display ("T=%0t [Generator] Wait for driver to be done", $time);
        @(drv_done);
        end
    endtask
    endclass


    // Lets say that the environment class was already there, and generator is 
    // a new component that needs to be included in the ENV. So a child ENV can
    // be derived and generator be instantiated in it along with all others.
    // Note that the run task should be overridden to start the generator as 
    // well.
    class env_w_gen extends env;
    generator g0;

    event drv_done;
    mailbox drv_mbx;

    function new();
        super.new();
        g0 = new;
        drv_mbx = new;
    endfunction

    virtual task run();
        // Connect virtual interface handles
        d0.vif = vif;
        m0.vif = vif;
        
        // Connect mailboxes between each component
        d0.drv_mbx = drv_mbx;
        g0.drv_mbx = drv_mbx;
        
        m0.scb_mbx = scb_mbx;
        s0.scb_mbx = scb_mbx;
        
        // Connect event handles
        d0.drv_done = drv_done;
        g0.drv_done = drv_done;
        
        // Start all components - a fork join_any is used because 
        // the stimulus is generated by the generator and we want the
        // simulation to exit only when the generator has finished 
        // creating all transactions. Until then all other components
        // have to run in the background.
        fork
            s0.run();
            d0.run();
            m0.run();
        g0.run();
        join_any
    endtask
endclass